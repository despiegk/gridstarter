module main

import os.cmdline
// import os
import freeflowuniverse.crystallib.actionrunner
import os

fn do() ! {

}

fn main() {
	do() or { panic(err) }
}
