module renumeration


struct Simulator{

}

struct Simulation{
	nr_people u32
	avg_monthly_points u8
	
}

pub fn (mut sim Simulator) calc(){
	
}