module postgresql

import freeflowuniverse.baobab.appsbox

// pub fn run( mut app appsbox.App)! {

// 	if app.wish == .build && app.build_state == .init {
// 		build(mut app)!
// 	}

// }

