module postgresql

