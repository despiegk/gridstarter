module appsbox

// import freeflowuniverse.crystallib.actionrunner
import freeflowuniverse.crystallib.pathlib
import regex

pub fn run (path0 string)!{

	mut path := pathlib.get_dir(path0, false)!	

	mut re := regex.regex_opt(".*") or {panic(err)}
	ar:=path.list(mut regex:re, 	recursive:true)!
	for p in ar{
		if p.path.ends_with(".md"){
			println(p)
		}
	}


}

// // set home directory and do initialization of multiple parts
// fn (mut apps AppsBox) home_set(path_ string) {
// 	mut path := path_
// 	if path == '' {
// 		// path="~/hub3"
// 		path = rootpath.rootdir()
// 	}
// 	if apps.apps_path == '' {
// 		apps.apps_path = path
// 	}
// 	if apps.bin_path == '' {
// 		apps.bin_path = '$apps.apps_path/bin'
// 	}
// 	if apps.var_path == '' {
// 		apps.var_path = '$apps.apps_path/var'
// 	}
// 	apps.apps_path = apps.apps_path.replace('~', os.home_dir())
// 	if !os.exists(apps.apps_path) {
// 		os.mkdir_all(apps.apps_path) or { panic('cannot create apps_path') }
// 	}
// 	apps.bin_path = apps.bin_path.replace('~', os.home_dir())
// 	if !os.exists(apps.bin_path) {
// 		os.mkdir_all(apps.bin_path) or { panic('cannot create bin_path') }
// 	}
// 	apps.var_path = apps.var_path.replace('~', os.home_dir())
// 	if !os.exists(apps.var_path) {
// 		os.mkdir_all(apps.var_path) or { panic('cannot create var_path') }
// 	}
// }
