module renumeration



