module appsbox


// import freeflowuniverse.crystallib.gridstarter.postgresql

// type MyApp = postgresql.
